library verilog;
use verilog.vl_types.all;
entity GATES_TT_vlg_vec_tst is
end GATES_TT_vlg_vec_tst;
